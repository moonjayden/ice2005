`timescale 1ns/1ns

module tb_custom;
	//clock
	reg CLK;
///////////////////////////////////////////////////
	//////////////////////////////////
	//Custom Module
	//input
	reg [7:0] a11, a12, a13, a14,
		  a21, a22, a23, a24,
		  a31, a32, a33, a34,
		  a41, a42, a43, a44;

    	reg [7:0] b11, b12, b13,
		  b21, b22, b23,
		  b31, b32, b33;

    	reg [3:0] S0_11, S0_12, S0_13,
   		  S0_21, S0_22, S0_23,
    		  S0_31, S0_32, S0_33;
	
	reg INIT;
	reg RST;
	reg PRESET;
	//output
	wire [7:0]OUT;
///////////////////////////////////////////////////
	//Module instantiation
	//Custom Module
	custom_module custom(
    	.a11(a11), .a12(a12), .a13(a13), .a14(a14),
    	.a21(a21), .a22(a22), .a23(a23), .a24(a24),
    	.a31(a31), .a32(a32), .a33(a33), .a34(a34),
    	.a41(a41), .a42(a42), .a43(a43), .a44(a44),
    	.b11(b11), .b12(b12), .b13(b13),
    	.b21(b21), .b22(b22), .b23(b23),
    	.b31(b31), .b32(b32), .b33(b33),
    	.clk(CLK), .init(INIT),
	.rst(RST), .preset(PRESET),
	.s0_11(S0_11), .s0_12(S0_12), .s0_13(S0_13),
    	.s0_21(S0_21), .s0_22(S0_22), .s0_23(S0_23),
    	.s0_31(S0_31), .s0_32(S0_32), .s0_33(S0_33),
    	.out(OUT));


///////////////////////////////////////////////////

	initial
	begin
		INIT = 1'b0;
    		RST = 1'b1;
    		PRESET = 1'b0;
    		CLK = 1'b0;
    		S0_11 = 4'b0000; S0_12 = 4'b0000; S0_13 = 4'b0000;
   		S0_21 = 4'b0000; S0_22 = 4'b0000; S0_23 = 4'b0000;
    		S0_31 = 4'b0000; S0_32 = 4'b0000; S0_33 = 4'b0000;

    		a11 = 8'd1; a12 = 8'd2; a13 = 8'd3; a14 = 8'd4;
		a21 = 8'd2; a22 = 8'd3; a23 = 8'd4; a24 = 8'd5;
		a31 = 8'd3; a32 = 8'd4; a33 = 8'd5; a34 = 8'd5;
		a41 = 8'd3; a42 = 8'd4; a43 = 8'd5; a44 = 8'd5;

		b11 = 8'd9; b12 = 8'd8; b13 = 8'd7;
		b21 = 8'd8; b22 = 8'd7; b23 = 8'd6;
		b31 = 8'd7; b32 = 8'd6; b33 = 8'd5;
		
		
	end

///////////////////////////////////////////////////  
	//Clock Cycle Time <- 20ns = 50MHz
	initial begin
    		forever begin
        		#10 CLK = ~CLK;
    		end
	end 		
///////////////////////////////////////////////////
	//test patterns
	initial 
	begin	
	//c11
		#20 RST = 1'b0;
    		 	S0_11 = 4'b0000; S0_12 = 4'b0100; S0_13 = 4'b1000;
   			S0_21 = 4'b0001; S0_22 = 4'b0101; S0_23 = 4'b1001;
    			S0_31 = 4'b0010; S0_32 = 4'b0110; S0_33 = 4'b1010;
		#20 INIT = 1'b1;
	//c12
		#20 INIT = 1'b0;
		 	S0_11 = 4'b0100; S0_12 = 4'b1000; S0_13 = 4'b1100;
   			S0_21 = 4'b0101; S0_22 = 4'b1001; S0_23 = 4'b1101;
    			S0_31 = 4'b0110; S0_32 = 4'b1010; S0_33 = 4'b1110;
    		#40 INIT = 1'b1;
		
	//c21
    		#20 INIT = 1'b0;
		 	S0_11 = 4'b0001; S0_12 = 4'b0101; S0_13 = 4'b1001;
   			S0_21 = 4'b0010; S0_22 = 4'b0110; S0_23 = 4'b1010;
    			S0_31 = 4'b0011; S0_32 = 4'b0111; S0_33 = 4'b1011;
		#20 INIT = 1'b1;
		
	//c22
    		#20 INIT = 1'b0; 
		 	S0_11 = 4'b0101; S0_12 = 4'b1001; S0_13 = 4'b1101;
   			S0_21 = 4'b0110; S0_22 = 4'b1010; S0_23 = 4'b1110;
    			S0_31 = 4'b0111; S0_32 = 4'b1011; S0_33 = 4'b1111;
    		#20 INIT = 1'b1;
		
	end
///////////////////////////////////////////////////
///////////////////////////////////////////////////////////////


endmodule
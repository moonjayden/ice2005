`timescale 1ns/1ns

module tb_parallel;
   //clock
   reg CLK;
///////////////////////////////////////////////////
   //////////////////////////////////
   //Custom Module
   //input
   //input
   reg [7:0] a11, a12, a13, a14,
        a21, a22, a23, a24,
        a31, a32, a33, a34,
        a41, a42, a43, a44;

       reg [7:0] b11, b12, b13,
        b21, b22, b23,
        b31, b32, b33;

       reg [3:0] S0, S1;
   reg WE_1, WE_2;
   reg RST;
   reg PRESET;
   //output
   wire [7:0]OUT;
///////////////////////////////////////////////////
   //Module instantiation
   //Custom Module
   Parallel_module parallel(
       .a11(a11), .a12(a12), .a13(a13), .a14(a14),
       .a21(a21), .a22(a22), .a23(a23), .a24(a24),
       .a31(a31), .a32(a32), .a33(a33), .a34(a34),
       .a41(a41), .a42(a42), .a43(a43), .a44(a44),
       .b11(b11), .b12(b12), .b13(b13),
       .b21(b21), .b22(b22), .b23(b23),
       .b31(b31), .b32(b32), .b33(b33),
   .s0(S0), .s1(S1),
       .clk(CLK), .we_1(WE_1), .we_2(WE_2),
   .rst(RST), .preset(PRESET),
       .out(OUT));


///////////////////////////////////////////////////

   initial
   begin
          RST = 1'b1;
          PRESET = 1'b0;
          CLK = 1'b0;
      WE_1=1'b0; WE_2=1'b0;
          //S0 = 4'b0000;
          S1 = 4'b0000;


          a11 = 8'd1; a12 = 8'd2; a13 = 8'd3; a14 = 8'd4;
      a21 = 8'd2; a22 = 8'd3; a23 = 8'd4; a24 = 8'd5;
      a31 = 8'd3; a32 = 8'd4; a33 = 8'd5; a34 = 8'd5;
      a41 = 8'd3; a42 = 8'd4; a43 = 8'd5; a44 = 8'd5;

      b11 = 8'd9; b12 = 8'd8; b13 = 8'd7;
      b21 = 8'd8; b22 = 8'd7; b23 = 8'd6;
      b31 = 8'd7; b32 = 8'd6; b33 = 8'd5;
      
      
   end

///////////////////////////////////////////////////  
   //Clock Cycle Time <- 20ns = 50MHz
   initial begin
          forever begin
              #10 CLK = ~CLK;
          end
   end       
///////////////////////////////////////////////////
   //test patterns
   initial 
   begin   
   //s0: 0->1->2->4->5->6->1->2->3->5->6->7->7->7->...->...
      #20 RST = 1'b0;
      #20 S1 = 4'b0010;
      #20 S1 = 4'b0001; WE_1=1'b1;
	#20 S1 = 4'b0000;
	#20 WE_1=1'b0; WE_2=1'b1;
          #20 S0 = 4'b0000; WE_2=1'b0;
          #20 S0 = 4'b0001;
          #20 S0 = 4'b0010;
          #20 S0 = 4'b0100;
          #20 S0 = 4'b0101;
          #20 S0 = 4'b0110;
          #20 S0 = 4'b0001;
          #20 S0 = 4'b0010;
      #20 S0 = 4'b0011;
          #20 S0 = 4'b0101;
          #20 S0 = 4'b0110;
          #20 S0 = 4'b0111;
   end
///////////////////////////////////////////////////
///////////////////////////////////////////////////////////////


endmodule
`timescale 1ns/1ns

module tb_pe_input;
	integer count;
	//clock
	reg CLK;
///////////////////////////////////////////////////
	//////////////////////////////////
	//input
	reg [7:0] a11, a12, a13, a14,
		  a21, a22, a23, a24,
		  a31, a32, a33, a34,
		  a41, a42, a43, a44;

    	reg [7:0] b11, b12, b13,
		  b21, b22, b23,
		  b31, b32, b33;

    	reg [3:0] S0, S1;
	
	
	//output
	wire [7:0] A_OUT, B_OUT;
	//////////////////////////////////

///////////////////////////////////////////////////
	//Module instantiation
	//PE Input Module
	pe_input_module pe_input(
	.a11(a11), .a12(a12), .a13(a13), .a14(a14),
    	.a21(a21), .a22(a22), .a23(a23), .a24(a24),
    	.a31(a31), .a32(a32), .a33(a33), .a34(a34),
    	.a41(a41), .a42(a42), .a43(a43), .a44(a44),
    	.b11(b11), .b12(b12), .b13(b13),
    	.b21(b21), .b22(b22), .b23(b23),
    	.b31(b31), .b32(b32), .b33(b33),
	.s0(S0), .s1(S1), .a_out(A_OUT), .b_out(B_OUT));
	

///////////////////////////////////////////////////
	initial
	begin
    		CLK = 1'b0;
    		a11 = 8'd1; a12 = 8'd2; a13 = 8'd3; a14 = 8'd4;
		a21 = 8'd2; a22 = 8'd3; a23 = 8'd4; a24 = 8'd5;
		a31 = 8'd3; a32 = 8'd4; a33 = 8'd5; a34 = 8'd5;
		a41 = 8'd3; a42 = 8'd4; a43 = 8'd5; a44 = 8'd5;

		b11 = 8'd9; b12 = 8'd8; b13 = 8'd7;
		b21 = 8'd8; b22 = 8'd7; b23 = 8'd6;
		b31 = 8'd7; b32 = 8'd6; b33 = 8'd5;

		S0 = 4'd0; S1 = 4'd0;

	end
///////////////////////////////////////////////////
	//Clock Cycle Time <- 20ns = 50MHz
	initial begin
    		forever begin
        		#10 CLK = ~CLK;
    		end
	end
///////////////////////////////////////////////////
	//Test Pattern
	initial
	begin
		#10;
		for (count = 0;count < 16;count=count+1)
		begin
			S0 <= count;
			S1 <= count;
			#10; 
		end
		#20 S0 = 4'b0100; S1 = 4'b0001;
    		#20 S0 = 4'b1000; S1 = 4'b0010;
    		#20 S0 = 4'b0001; S1 = 4'b0100;
    		#20 S0 = 4'b0101; S1 = 4'b0101;
    		#20 S0 = 4'b1001; S1 = 4'b0110;
    		#20 S0 = 4'b0010; S1 = 4'b1000;
    		#20 S0 = 4'b0110; S1 = 4'b1001;
    		#20 S0 = 4'b1010; S1 = 4'b1010;

	end
///////////////////////////////////////////////////

	
endmodule
